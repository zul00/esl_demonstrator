LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY PulseWidthModulator IS
  PORT (
         pulse : OUT std_logic;
         clk : IN std_logic
       );
END ENTITY;

ARCHITECTURE bhv OF PulseWidthModulator IS
BEGIN
END ARCHITECTURE bhv;
